netcdf lfric_xios_write_test {
dimensions:
	axis_nbounds = 2 ;
	Two = 2 ;
	nMesh2d_node = 1 ;
	nMesh2d_edge = UNLIMITED ; // (0 currently)
	nMesh2d_face = 9 ;
	nMesh2d_vertex = 4 ;
	vert_axis_half_levels = 5 ;
	time = UNLIMITED ; // (10 currently)
variables:
	int Mesh2d ;
		Mesh2d:cf_role = "mesh_topology" ;
		Mesh2d:long_name = "Topology data of 2D unstructured mesh" ;
		Mesh2d:topology_dimension = 2 ;
		Mesh2d:node_coordinates = "Mesh2d_node_x Mesh2d_node_y" ;
		Mesh2d:edge_coordinates = "Mesh2d_edge_x Mesh2d_edge_y" ;
		Mesh2d:edge_node_connectivity = "Mesh2d_edge_nodes" ;
		Mesh2d:face_edge_connectivity = "Mesh2d_face_edges" ;
		Mesh2d:edge_face_connectivity = "Mesh2d_edge_face_links" ;
		Mesh2d:face_face_connectivity = "Mesh2d_face_links" ;
		Mesh2d:face_coordinates = "Mesh2d_face_x Mesh2d_face_y" ;
		Mesh2d:face_node_connectivity = "Mesh2d_face_nodes" ;
		Mesh2d:geometry = "planar" ;
	float Mesh2d_node_x(nMesh2d_node) ;
		Mesh2d_node_x:standard_name = "projection_x_coordinate" ;
		Mesh2d_node_x:long_name = "x coordinate of projection" ;
		Mesh2d_node_x:units = "m" ;
		Mesh2d_node_x:scale_factor = 10000. ;
	float Mesh2d_node_y(nMesh2d_node) ;
		Mesh2d_node_y:standard_name = "projection_y_coordinate" ;
		Mesh2d_node_y:long_name = "y coordinate of projection" ;
		Mesh2d_node_y:units = "m" ;
		Mesh2d_node_y:scale_factor = 10000. ;
	float Mesh2d_edge_x(nMesh2d_edge) ;
		Mesh2d_edge_x:standard_name = "projection_x_coordinate" ;
		Mesh2d_edge_x:long_name = "x coordinate of projection" ;
		Mesh2d_edge_x:units = "m" ;
		Mesh2d_edge_x:scale_factor = 10000. ;
	float Mesh2d_edge_y(nMesh2d_edge) ;
		Mesh2d_edge_y:standard_name = "projection_y_coordinate" ;
		Mesh2d_edge_y:long_name = "y coordinate of projection" ;
		Mesh2d_edge_y:units = "m" ;
		Mesh2d_edge_y:scale_factor = 10000. ;
	int Mesh2d_edge_nodes(nMesh2d_edge, Two) ;
		Mesh2d_edge_nodes:cf_role = "edge_node_connectivity" ;
		Mesh2d_edge_nodes:long_name = "Maps every edge/link to two nodes that it connects." ;
		Mesh2d_edge_nodes:start_index = 0 ;
	float Mesh2d_face_x(nMesh2d_face) ;
		Mesh2d_face_x:standard_name = "projection_x_coordinate" ;
		Mesh2d_face_x:long_name = "x coordinate of projection" ;
		Mesh2d_face_x:units = "m" ;
		Mesh2d_face_x:scale_factor = 10000. ;
	float Mesh2d_face_y(nMesh2d_face) ;
		Mesh2d_face_y:standard_name = "projection_y_coordinate" ;
		Mesh2d_face_y:long_name = "y coordinate of projection" ;
		Mesh2d_face_y:units = "m" ;
		Mesh2d_face_y:scale_factor = 10000. ;
	int Mesh2d_face_nodes(nMesh2d_face, nMesh2d_vertex) ;
		Mesh2d_face_nodes:cf_role = "face_node_connectivity" ;
		Mesh2d_face_nodes:long_name = "Maps every face to its corner nodes." ;
		Mesh2d_face_nodes:start_index = 0 ;
	int Mesh2d_face_edges(nMesh2d_face, nMesh2d_vertex) ;
		Mesh2d_face_edges:cf_role = "face_edge_connectivity" ;
		Mesh2d_face_edges:long_name = "Maps every face to its edges." ;
		Mesh2d_face_edges:start_index = 0 ;
		Mesh2d_face_edges:_FillValue = 999999 ;
	int Mesh2d_edge_face_links(nMesh2d_edge, Two) ;
		Mesh2d_edge_face_links:cf_role = "edge_face_connectivity" ;
		Mesh2d_edge_face_links:long_name = "neighbor faces for edges" ;
		Mesh2d_edge_face_links:start_index = 0 ;
		Mesh2d_edge_face_links:_FillValue = -999 ;
		Mesh2d_edge_face_links:comment = "missing neighbor faces are indicated using _FillValue" ;
	int Mesh2d_face_links(nMesh2d_face, nMesh2d_vertex) ;
		Mesh2d_face_links:cf_role = "face_face_connectivity" ;
		Mesh2d_face_links:long_name = "Indicates which other faces neighbor each face" ;
		Mesh2d_face_links:start_index = 0 ;
		Mesh2d_face_links:_FillValue = 999999 ;
		Mesh2d_face_links:flag_values = -1 ;
		Mesh2d_face_links:flag_meanings = "out_of_mesh" ;
	float vert_axis_half_levels(vert_axis_half_levels) ;
		vert_axis_half_levels:name = "vert_axis_half_levels" ;
	double time(time) ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:long_name = "Time axis" ;
		time:calendar = "gregorian" ;
		time:units = "seconds since 2024-01-01 15:00:00" ;
		time:time_origin = "2024-01-01 15:00:00" ;
		time:bounds = "time_bounds" ;
		time:coordinates = " forecast_reference_time forecast_period" ;
	double time_bounds(time, axis_nbounds) ;
		time_bounds:coordinates = " forecast_reference_time forecast_period" ;
	double temporal_field(time, vert_axis_half_levels, nMesh2d_face) ;
		temporal_field:mesh = "Mesh2d" ;
		temporal_field:location = "face" ;
		temporal_field:online_operation = "instant" ;
		temporal_field:interval_operation = "60 s" ;
		temporal_field:interval_write = "60 s" ;
		temporal_field:cell_methods = "time: point" ;
		temporal_field:coordinates = "Mesh2d_face_y Mesh2d_face_x forecast_reference_time forecast_period" ;
	double forecast_reference_time ;
		forecast_reference_time:units = "seconds since 2024-01-01 15:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
	double forecast_period(time) ;
		forecast_period:units = "seconds" ;
		forecast_period:standard_name = "forecast_period" ;
		forecast_period:coordinates = " forecast_reference_time forecast_period" ;

// global attributes:
		:name = "lfric_xios_write_test" ;
		:title = "Created by xios" ;
		:timeStamp = "2025-Feb-26 11:47:23 GMT" ;
		:uuid = "4f0f6d47-9240-4356-b1f6-b02f8adc4fe4" ;
		:description = "LFRic file format v0.2.0" ;
		:Conventions = "UGRID-1.0" ;
data:

 Mesh2d = 13795354 ;

 Mesh2d_node_x = 0 ;

 Mesh2d_node_y = 0 ;

 Mesh2d_face_x = 0.0001, 0.0002, 0.0001, 0.0003, 0.0001, 0.0003, 0.0002, 
    0.0003, 0.0002 ;

 Mesh2d_face_y = 0.0001, 0.0001, 0.0001, 0.0002, 0.0002, 0.0002, 0.0003, 
    0.0003, 0.0003 ;

 Mesh2d_face_nodes =
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;

 Mesh2d_face_edges =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 Mesh2d_face_links =
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _,
  _, _, _, _ ;

 vert_axis_half_levels = 0.5, 1.5, 2.5, 3.5, 4.5 ;

 time = 60, 120, 180, 240, 300, 360, 420, 480, 540, 600 ;

 time_bounds =
  60, 60,
  120, 120,
  180, 180,
  240, 240,
  300, 300,
  360, 360,
  420, 420,
  480, 480,
  540, 540,
  600, 600 ;

 temporal_field =
  20, 20, 20, 20, 20, 20, 20, 20, 20,
  20, 20, 20, 20, 20, 20, 20, 20, 20,
  20, 20, 20, 20, 20, 20, 20, 20, 20,
  20, 20, 20, 20, 20, 20, 20, 20, 20,
  20, 20, 20, 20, 20, 20, 20, 20, 20,
  6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667,
  6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667,
  6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667,
  6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667,
  6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667, 6.66666666666667, 6.66666666666667, 6.66666666666667, 
    6.66666666666667,
  26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667,
  26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667,
  26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667,
  26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667,
  26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667, 26.6666666666667, 26.6666666666667, 26.6666666666667, 
    26.6666666666667,
  5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333,
  5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333,
  5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333,
  5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333,
  5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333, 5.33333333333333, 5.33333333333333, 5.33333333333333, 
    5.33333333333333,
  32, 32, 32, 32, 32, 32, 32, 32, 32,
  32, 32, 32, 32, 32, 32, 32, 32, 32,
  32, 32, 32, 32, 32, 32, 32, 32, 32,
  32, 32, 32, 32, 32, 32, 32, 32, 32,
  32, 32, 32, 32, 32, 32, 32, 32, 32,
  4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857,
  4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857,
  4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857,
  4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857,
  4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857, 4.57142857142857, 4.57142857142857, 4.57142857142857, 
    4.57142857142857,
  36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286,
  36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286,
  36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286,
  36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286,
  36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286, 36.5714285714286, 36.5714285714286, 36.5714285714286, 
    36.5714285714286,
  4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206,
  4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206,
  4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206,
  4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206,
  4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206, 4.06349206349206, 4.06349206349206, 4.06349206349206, 
    4.06349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 0,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206,
  40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206, 40.6349206349206, 40.6349206349206, 40.6349206349206, 
    40.6349206349206 ;

 forecast_reference_time = 0 ;

 forecast_period = 60, 120, 180, 240, 300, 360, 420, 480, 540, 600 ;
}
